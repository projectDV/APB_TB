package apb_pkg;
`include "apn_txn"
`include "apb_gen"
`include "apb_drv"
`include "apb_mon"
`include "apb_txn"
`include "apb_rm"
`include "apb_sb"
`include "apb_env"
endpackage
